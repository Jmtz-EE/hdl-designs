module not_4 (
    input[3:0] a,b,
    output[3:0] x,y
);
    assign x = ~a;
    assign y = ~b; 
endmodule